BZh91AY&SY�+�  �_�Py��g߰����PX�w�anA(SH��OL"z���C@ dC�=@��$z���~��     " ��<��i=Q�� 4d40&&�	�&L�&	����CI�2h'�d�A�h �@h�+߈�*
������+��blI��С"ƒ�j�*�c\;��8'Dl�
h��WԺ�>�xv��n7d��]�;�%��F��&r�P���9$�-���41)F<GKu���ȿ�u�F�������Õ�#߾C�8���j�����M{�AƱci�� gVӑ�?�c�+�3�$��O\���u=���ƎI &�D8x���$��GpF�1�Y)w��P�N_�G[vzF%���V���c���q�.M~Nr�(��c.��Sa�/֛�2��� �EV%K��T��ru5����Bj�1�&ܶ*�`B���� b�@�p?6 ,$7��
��0��4R5aa�<�׾�NW�	q�%4�8�Lm���S�Mmu�H2���xo&�/QJ�!��)F'�v|��$yJ���)��pe�@,��,(ٝR`���f� ��D��I�d���-{=)0*be���L&?��踜���f:3�i�0[W0�nV-. 4V�hA��\#��<�I�c!l�pf���
��%*'i6@����V1d��r�:&n�x�[1��u���%E�c5�G=��Rg���!$�I5=/Z���+*�1���X�*��ƪ��Je�@L�().�p���D���+}��,�Ɉ�Z�!�t�&�aSh��}d4��.�x����s�fQK#�X8�2�ce���~Bx��Ľ��d}!���{�f�K �](��.�p�!<WN